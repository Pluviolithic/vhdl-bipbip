library IEEE;
use IEEE.numeric_bit.all;

entity s_box is
    port (
        x : in bit_vector(5 downto 0);
        y_out : out bit_vector(5 downto 0)
    );
end s_box;

-- change this to operate from memory
architecture lut of s_box is
    signal y : bit_vector(5 downto 0);
begin
    process (x) is
    begin
        case x is
            when "000000" => y <= "000000";
            when "000001" => y <= "000001";
            when "000010" => y <= "000010";
            when "000011" => y <= "000011";
            when "000100" => y <= "000100";
            when "000101" => y <= "000110";
            when "000110" => y <= "111110";
            when "000111" => y <= "111100";
            when "001000" => y <= "001000";
            when "001001" => y <= "010001";
            when "001010" => y <= "001110";
            when "001011" => y <= "010111";
            when "001100" => y <= "101011";
            when "001101" => y <= "110011";
            when "001110" => y <= "110101";
            when "001111" => y <= "101101";
            when "010000" => y <= "011001";
            when "010001" => y <= "011100";
            when "010010" => y <= "001001";
            when "010011" => y <= "001100";
            when "010100" => y <= "010101";
            when "010101" => y <= "010011";
            when "010110" => y <= "111101";
            when "010111" => y <= "111011";
            when "011000" => y <= "110001";
            when "011001" => y <= "101100";
            when "011010" => y <= "100101";
            when "011011" => y <= "111000";
            when "011100" => y <= "111010";
            when "011101" => y <= "100110";
            when "011110" => y <= "110110";
            when "011111" => y <= "101010";
            when "100000" => y <= "110100";
            when "100001" => y <= "011101";
            when "100010" => y <= "110111";
            when "100011" => y <= "011110";
            when "100100" => y <= "110000";
            when "100101" => y <= "011010";
            when "100110" => y <= "001011";
            when "100111" => y <= "100001";
            when "101000" => y <= "101110";
            when "101001" => y <= "011111";
            when "101010" => y <= "101001";
            when "101011" => y <= "011000";
            when "101100" => y <= "001111";
            when "101101" => y <= "111111";
            when "101110" => y <= "010000";
            when "101111" => y <= "100000";
            when "110000" => y <= "101000";
            when "110001" => y <= "000101";
            when "110010" => y <= "111001";
            when "110011" => y <= "010100";
            when "110100" => y <= "100100";
            when "110101" => y <= "001010";
            when "110110" => y <= "001101";
            when "110111" => y <= "100011";
            when "111000" => y <= "010010";
            when "111001" => y <= "100111";
            when "111010" => y <= "000111";
            when "111011" => y <= "110010";
            when "111100" => y <= "011011";
            when "111101" => y <= "101111";
            when "111110" => y <= "010110";
            when "111111" => y <= "100010";
        end case;
    end process;
    y_out <= y;
end lut;