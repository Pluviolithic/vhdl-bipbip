library IEEE;
use IEEE.numeric_bit.all;

entity pi_5 is
    port (
        x : in bit_vector(52 downto 0);
        y : out bit_vector(52 downto 0)
    );
end pi_5;

architecture Behavioral of pi_5 is
begin
    y(0) <= x(0);
    y(1) <= x(11);
    y(2) <= x(22);
    y(3) <= x(33);
    y(4) <= x(44);
    y(5) <= x(0);
    y(6) <= x(11);
    y(7) <= x(22);
    y(8) <= x(33);
    y(9) <= x(44);
    y(10) <= x(0);
    y(11) <= x(11);
    y(12) <= x(22);
    y(13) <= x(33);
    y(14) <= x(44);
    y(15) <= x(0);
    y(16) <= x(11);
    y(17) <= x(22);
    y(18) <= x(33);
    y(19) <= x(44);
    y(20) <= x(0);
    y(21) <= x(11);
    y(22) <= x(22);
    y(23) <= x(33);
    y(24) <= x(44);
    y(25) <= x(0);
    y(26) <= x(11);
    y(27) <= x(22);
    y(28) <= x(33);
    y(29) <= x(44);
    y(30) <= x(0);
    y(31) <= x(11);
    y(32) <= x(22);
    y(33) <= x(33);
    y(34) <= x(44);
    y(35) <= x(0);
    y(36) <= x(11);
    y(37) <= x(22);
    y(38) <= x(33);
    y(39) <= x(44);
    y(40) <= x(0);
    y(41) <= x(11);
    y(42) <= x(22);
    y(43) <= x(33);
    y(44) <= x(44);
    y(45) <= x(0);
    y(46) <= x(11);
    y(47) <= x(22);
    y(48) <= x(33);
    y(49) <= x(44);
    y(50) <= x(0);
    y(51) <= x(11);
    y(52) <= x(22);
end Behavioral;